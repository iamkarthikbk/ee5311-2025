** sch_path: /home/ee24s053/ee5311-2025/tut6/incr/step4_again/fa.sch
.subckt fa a b cin DGND DVDD cout_n
*.PININFO a:I b:I cin:I DGND:B DVDD:B cout_n:O
XM15 cout_n cin net1 DVDD sky130_fd_pr__pfet_01v8 L=0.15 W=1.68 nf=1 m=1
XM16 net1 b DVDD DVDD sky130_fd_pr__pfet_01v8 L=0.15 W=3.36 nf=1 m=1
XM17 net1 a DVDD DVDD sky130_fd_pr__pfet_01v8 L=0.15 W=3.36 nf=1 m=1
XM18 cout_n cin net2 DGND sky130_fd_pr__nfet_01v8 L=0.15 W=0.84 nf=1 m=1
XM19 net2 b DGND DGND sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM20 net2 a DGND DGND sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM21 net4 a DVDD DVDD sky130_fd_pr__pfet_01v8 L=0.15 W=1.68 nf=1 m=1
XM22 cout_n b net4 DVDD sky130_fd_pr__pfet_01v8 L=0.15 W=1.68 nf=1 m=1
XM23 cout_n b net3 DGND sky130_fd_pr__nfet_01v8 L=0.15 W=0.84 nf=1 m=1
XM24 net3 a DGND DGND sky130_fd_pr__nfet_01v8 L=0.15 W=0.84 nf=1 m=1
.ends
.end
