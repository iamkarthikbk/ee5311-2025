** sch_path: /home/ee24s053/ee5311-2025/tut6/rca/rca8b_tb.sch
**.subckt rca8b_tb
x1 GND GND GND GND GND GND GND GND VDD VDD VDD VDD VDD VDD VDD VDD VDD cout_tap cin_tap GND s7_tap net1 net2 net3 net4 net5 net6
+ net7 rca8b
V1 cin_tap GND PULSE(0 1.8 0 5ps 5ps 1ns 2ns)
V2 VDD GND 1.8
x2 VDD cout_tap net8 GND invx1
x3 VDD s7_tap net9 GND invx1
**** begin user architecture code
.lib /cad/share/pdk/sky130B/libs.tech/combined/sky130.lib.spice tt


.include /home/ee24s053/ee5311-2025/tut6/rca/rca8b_extracted.spice
.control
tran 1p 20n
plot v(s7_tap) v(cout_tap)
meas tran tlh_carry trig v(cin_tap) val=0.9 rise=1 targ v(cout_tap) val=0.9 rise=1
meas tran thl_carry trig v(cin_tap) val=0.9 fall=1 targ v(cout_tap) val=0.9 fall=1
let carry_delay = ($&tlh_carry + $&thl_carry)/2
echo carry delay: $&carry_delay
meas tran tlh_sum trig v(cin_tap) val=0.9 rise=1 targ v(s7_tap) val=0.9 rise=1
meas tran thl_sum trig v(cin_tap) val=0.9 fall=1 targ v(s7_tap) val=0.9 fall=1
let sum_delay = ($&tlh_sum + $&thl_sum)/2
echo sum delay: $&sum_delay
.endc

**** end user architecture code
**.ends

* expanding   symbol:  /home/ee24s053/ee5311-2025/tut6/again/inv/invx1.sym # of pins=4
** sym_path: /home/ee24s053/ee5311-2025/tut6/again/inv/invx1.sym
** sch_path: /home/ee24s053/ee5311-2025/tut6/again/inv/invx1.sch
.subckt invx1 DVDD in out DGND
*.ipin in
*.opin out
*.iopin DVDD
*.iopin DGND
XM2 out in DVDD DVDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.84 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM1 out in DGND DGND sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends

.GLOBAL VDD
.GLOBAL GND
.end
