** sch_path: /home/ee24s053/ee5311-2025/tut1/tut1-expt3.sch
**.subckt tut1-expt3
Vin1 Vin GND 1.8
Vdd1 net1 GND 1.8
XM1 net1 Vin GND GND sky130_fd_pr__nfet_01v8 L={Length} W={Width} nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
**** begin user architecture code
.lib /cad/share/pdk/sky130B/libs.tech/combined/sky130.lib.spice tt


.param Width = 0.42
.param Length = 0.15
.dc Vdd1 0 1.8 0.01
.control
  let index = 1
  set cache = ''
  while index <= 10
    let newW = index * 0.42
    let newL = index * 0.15
    alterparam Width = $&newW
    alterparam Length = $&newL
    reset
    run
    set cache = ( $cache dc{$&index}.i(VDD1)*-1 )
    let index = index + 1
end
plot $cache
.endc


**** end user architecture code
**.ends
.GLOBAL GND
.end
