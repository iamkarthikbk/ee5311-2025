* NGSPICE file created from nand2x1.ext - technology: sky130A
.subckt nand2x1 DVDD DGND A B F
X0 F.t3 A.t0 a_n694_n141# DGND.t1 sky130_fd_pr__nfet_01v8 ad=0.21 pd=1.34 as=0.252 ps=2.28 w=0.84 l=0.15
X1 a_n694_n141# A.t1 F.t2 DGND.t0 sky130_fd_pr__nfet_01v8 ad=0.252 pd=2.28 as=0.21 ps=1.34 w=0.84 l=0.15
X2 F.t1 A.t2 DVDD.t3 DVDD.t2 sky130_fd_pr__pfet_01v8 ad=0.21 pd=1.34 as=0.252 ps=2.28 w=0.84 l=0.15
X3 DVDD.t1 A.t3 F.t0 DVDD.t0 sky130_fd_pr__pfet_01v8 ad=0.5166 pd=2.07 as=0.21 ps=1.34 w=0.84 l=0.15
X4 a_n694_n141# B.t0 DGND.t5 DGND.t4 sky130_fd_pr__nfet_01v8 ad=0.21 pd=1.34 as=0.252 ps=2.28 w=0.84 l=0.15
X5 F.t5 B.t1 DVDD.t7 DVDD.t6 sky130_fd_pr__pfet_01v8 ad=0.21 pd=1.34 as=0.5166 ps=2.07 w=0.84 l=0.15
X6 DGND.t3 B.t2 a_n694_n141# DGND.t2 sky130_fd_pr__nfet_01v8 ad=0.252 pd=2.28 as=0.21 ps=1.34 w=0.84 l=0.15
X7 DVDD.t5 B.t3 F.t4 DVDD.t4 sky130_fd_pr__pfet_01v8 ad=0.252 pd=2.28 as=0.21 ps=1.34 w=0.84 l=0.15
R0 A.t3 A.t1 557.514
R1 A.t2 A.t3 526.987
R2 A.n0 A.t0 253.304
R3 A.n0 A.t2 251.697
R4 A A.n0 152.475
R5 F F.n0 400.771
R6 F.n3 F.n1 324.349
R7 F.n3 F.n2 164.321
R8 F F.n3 76.424
R9 F.n0 F.t4 58.6315
R10 F.n0 F.t5 58.6315
R11 F.n1 F.t0 58.6315
R12 F.n1 F.t1 58.6315
R13 F.n2 F.t2 35.7148
R14 F.n2 F.t3 35.7148
R15 DGND DGND.t2 4633.85
R16 DGND.t4 DGND.t0 3930.1
R17 DGND.t2 DGND.t4 1851.13
R18 DGND.t0 DGND.t1 1851.13
R19 DGND.n0 DGND.t5 165.412
R20 DGND.n0 DGND.t3 165.126
R21 DGND DGND.n0 0.251802
R22 DVDD DVDD.t4 945.405
R23 DVDD.t6 DVDD.t0 809.26
R24 DVDD.n1 DVDD.t3 405.666
R25 DVDD.n2 DVDD.t5 405.378
R26 DVDD.t4 DVDD.t6 381.173
R27 DVDD.t0 DVDD.t2 381.173
R28 DVDD.n1 DVDD.n0 346.253
R29 DVDD.n0 DVDD.t7 253.286
R30 DVDD.n0 DVDD.t1 35.1791
R31 DVDD.n2 DVDD.n1 0.529146
R32 DVDD DVDD.n2 0.2505
R33 B.t1 B.t0 557.514
R34 B.t3 B.t1 526.987
R35 B.n0 B.t2 253.304
R36 B.n0 B.t3 251.697
R37 B B.n0 152.388
C0 F A 0.074645f
C1 F DVDD 0.289908f
C2 a_n694_n141# A 0.047483f
C3 DVDD a_n694_n141# 0.048333f
C4 B F 0.03475f
C5 DVDD A 0.2002f
C6 B a_n694_n141# 0.028801f
C7 F a_n694_n141# 0.211072f
C8 B A 0.017336f
C9 B DVDD 0.207843f
C10 F DGND 0.134889f
C11 B DGND 0.350349f
C12 A DGND 0.320413f
C13 DVDD DGND 1.43629f
C14 a_n694_n141# DGND 0.495326f
.ends
