* NGSPICE file created from fa.ext - technology: sky130A

.subckt fa sum_n a cout_n b cin DVDD DGND
X0 a_n2273_210# cin cout_n DVDD sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X1 cout_n b a_n2493_n118# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.105 ps=0.92 w=0.42 l=0.15
X2 a_n2183_210# a a_n2273_210# DVDD sky130_fd_pr__pfet_01v8 ad=0.21 pd=1.34 as=0.126 ps=1.14 w=0.84 l=0.15
X3 a_81_210# a a_n49_210# DVDD sky130_fd_pr__pfet_01v8 ad=0.21 pd=1.34 as=0.21 ps=1.34 w=0.84 l=0.15
X4 a_n2053_n118# a a_n2183_n118# DGND sky130_fd_pr__nfet_01v8 ad=0.105 pd=0.92 as=0.105 ps=0.92 w=0.42 l=0.15
X5 a_n1573_n118# b a_n1703_n118# DGND sky130_fd_pr__nfet_01v8 ad=0.105 pd=0.92 as=0.105 ps=0.92 w=0.42 l=0.15
X6 a_n49_n118# a a_n139_n118# DGND sky130_fd_pr__nfet_01v8 ad=0.105 pd=0.92 as=0.063 ps=0.72 w=0.42 l=0.15
X7 a_n1109_210# cin DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.252 ps=2.28 w=0.84 l=0.15
X8 a_n1923_210# a a_n2053_210# DVDD sky130_fd_pr__pfet_01v8 ad=0.21 pd=1.34 as=0.21 ps=1.34 w=0.84 l=0.15
X9 a_n1443_210# b a_n1573_210# DVDD sky130_fd_pr__pfet_01v8 ad=0.21 pd=1.34 as=0.21 ps=1.34 w=0.84 l=0.15
X10 a_n669_210# a DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.21 ps=1.34 w=0.84 l=0.15
X11 DVDD b a_n1109_210# DVDD sky130_fd_pr__pfet_01v8 ad=0.21 pd=1.34 as=0.126 ps=1.14 w=0.84 l=0.15
X12 a_n269_n118# b a_n399_n118# DGND sky130_fd_pr__nfet_01v8 ad=0.105 pd=0.92 as=0.105 ps=0.92 w=0.42 l=0.15
X13 DVDD a a_n1923_210# DVDD sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.21 ps=1.34 w=0.84 l=0.15
X14 a_n2273_210# b a_n1443_210# DVDD sky130_fd_pr__pfet_01v8 ad=0.252 pd=2.28 as=0.21 ps=1.34 w=0.84 l=0.15
X15 a_n669_n118# a DGND DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.105 ps=0.92 w=0.42 l=0.15
X16 a_n1703_210# b DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.21 pd=1.34 as=0.126 ps=1.14 w=0.84 l=0.15
X17 a_n1109_210# b DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.21 ps=1.34 w=0.84 l=0.15
X18 a_n49_210# a a_n139_210# DVDD sky130_fd_pr__pfet_01v8 ad=0.21 pd=1.34 as=0.126 ps=1.14 w=0.84 l=0.15
X19 a_n139_n118# b a_n269_n118# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.105 ps=0.92 w=0.42 l=0.15
X20 a_n1573_210# b a_n1703_210# DVDD sky130_fd_pr__pfet_01v8 ad=0.21 pd=1.34 as=0.21 ps=1.34 w=0.84 l=0.15
X21 DVDD a a_n1109_210# DVDD sky130_fd_pr__pfet_01v8 ad=0.21 pd=1.34 as=0.126 ps=1.14 w=0.84 l=0.15
X22 a_n269_210# b a_n399_210# DVDD sky130_fd_pr__pfet_01v8 ad=0.21 pd=1.34 as=0.21 ps=1.34 w=0.84 l=0.15
X23 a_81_n118# a a_n49_n118# DGND sky130_fd_pr__nfet_01v8 ad=0.105 pd=0.92 as=0.105 ps=0.92 w=0.42 l=0.15
X24 a_n139_210# b a_n269_210# DVDD sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.21 ps=1.34 w=0.84 l=0.15
X25 sum_n cout_n a_n669_210# DVDD sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X26 a_n1443_n118# b a_n1573_n118# DGND sky130_fd_pr__nfet_01v8 ad=0.105 pd=0.92 as=0.105 ps=0.92 w=0.42 l=0.15
X27 a_n489_210# cin sum_n DVDD sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.126 ps=1.14 w=0.84 l=0.15
X28 a_n2713_n118# a DGND DGND sky130_fd_pr__nfet_01v8 ad=0.105 pd=0.92 as=0.126 ps=1.44 w=0.42 l=0.15
X29 a_n399_210# b a_n489_210# DVDD sky130_fd_pr__pfet_01v8 ad=0.21 pd=1.34 as=0.126 ps=1.14 w=0.84 l=0.15
X30 DVDD a a_81_210# DVDD sky130_fd_pr__pfet_01v8 ad=0.252 pd=2.28 as=0.21 ps=1.34 w=0.84 l=0.15
X31 a_n2273_n118# b a_n1443_n118# DGND sky130_fd_pr__nfet_01v8 ad=0.126 pd=1.44 as=0.105 ps=0.92 w=0.42 l=0.15
X32 a_n2493_n118# b a_n2583_n118# DGND sky130_fd_pr__nfet_01v8 ad=0.105 pd=0.92 as=0.063 ps=0.72 w=0.42 l=0.15
X33 DGND a a_81_n118# DGND sky130_fd_pr__nfet_01v8 ad=0.126 pd=1.44 as=0.105 ps=0.92 w=0.42 l=0.15
X34 a_n2183_n118# a a_n2273_n118# DGND sky130_fd_pr__nfet_01v8 ad=0.105 pd=0.92 as=0.063 ps=0.72 w=0.42 l=0.15
X35 cout_n b a_n2493_210# DVDD sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.21 ps=1.34 w=0.84 l=0.15
X36 a_n2583_n118# a a_n2713_n118# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.105 ps=0.92 w=0.42 l=0.15
X37 a_n2273_n118# cin cout_n DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X38 a_n2713_210# a DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.21 pd=1.34 as=0.252 ps=2.28 w=0.84 l=0.15
X39 DGND b a_n1109_n118# DGND sky130_fd_pr__nfet_01v8 ad=0.105 pd=0.92 as=0.063 ps=0.72 w=0.42 l=0.15
X40 a_n399_n118# b a_n489_n118# DGND sky130_fd_pr__nfet_01v8 ad=0.105 pd=0.92 as=0.063 ps=0.72 w=0.42 l=0.15
X41 DGND a a_n1109_n118# DGND sky130_fd_pr__nfet_01v8 ad=0.105 pd=0.92 as=0.063 ps=0.72 w=0.42 l=0.15
X42 a_n2583_210# a a_n2713_210# DVDD sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.21 ps=1.34 w=0.84 l=0.15
X43 a_n2053_210# a a_n2183_210# DVDD sky130_fd_pr__pfet_01v8 ad=0.21 pd=1.34 as=0.21 ps=1.34 w=0.84 l=0.15
X44 a_n1923_n118# a a_n2053_n118# DGND sky130_fd_pr__nfet_01v8 ad=0.105 pd=0.92 as=0.105 ps=0.92 w=0.42 l=0.15
X45 a_n1109_n118# cin DGND DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.126 ps=1.44 w=0.42 l=0.15
X46 a_n489_n118# cin sum_n DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X47 a_n2493_210# b a_n2583_210# DVDD sky130_fd_pr__pfet_01v8 ad=0.21 pd=1.34 as=0.126 ps=1.14 w=0.84 l=0.15
X48 a_n1109_n118# b DGND DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.105 ps=0.92 w=0.42 l=0.15
X49 sum_n cout_n a_n669_n118# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.063 ps=0.72 w=0.42 l=0.15
X50 a_n1703_n118# b DGND DGND sky130_fd_pr__nfet_01v8 ad=0.105 pd=0.92 as=0.063 ps=0.72 w=0.42 l=0.15
X51 DGND a a_n1923_n118# DGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.105 ps=0.92 w=0.42 l=0.15
.ends

