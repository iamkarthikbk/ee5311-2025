** sch_path: /home/ee24s053/ee5311-2025/tut4/expt2/ro9.sch
**.subckt ro9
x1 net1 vout inv
x2 net2 net1 inv
x3 net3 net2 inv
x4 net4 net3 inv
x5 net5 net4 inv
x6 net6 net5 inv
x7 net7 net6 inv
Vdd1 VDD GND {vdd_val}
x8 net8 net7 inv
x9 vout net8 inv
**** begin user architecture code
.lib /cad/share/pdk/sky130B/libs.tech/combined/sky130.lib.spice tt


.param wp = 0.84
.param vdd_val = 1.8
.ic v(vout) = 0
.control
let lv_iters = 9
let v_vdd = vector(lv_iters)
let v_period = vector(lv_iters)
let v_freq = vector(lv_iters)
let lv_index = 0
while lv_index < lv_iters
	let lv_vdd = 1.0 + (lv_index * 0.1)
	let vhalf = lv_vdd / 2
	alterparam vdd_val = $&lv_vdd
	reset
	tran 1p 10n
	meas tran prd trig v(vout) val=vhalf rise=3 targ v(vout) val=vhalf rise=4
	let v_period[lv_index] = $&prd
	let v_freq[lv_index] = 1/$&prd
	let v_vdd[lv_index] = $&lv_vdd
	let lv_index = lv_index + 1
end
plot v_period vs v_vdd
plot v_freq vs v_vdd
.endc


**** end user architecture code
**.ends

* expanding   symbol:  /home/ee24s053/ee5311-2025/tut3/syms/inv.sym # of pins=2
** sym_path: /home/ee24s053/ee5311-2025/tut3/syms/inv.sym
** sch_path: /home/ee24s053/ee5311-2025/tut3/syms/inv.sch
.subckt inv out in
*.ipin in
*.opin out
XM1 out in VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W={wp} nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 out in GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends

.GLOBAL VDD
.GLOBAL GND
.end
