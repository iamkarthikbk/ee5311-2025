** sch_path: /home/ee24s053/ee5311-2025/tut5/inv/prim/inv.sch
.subckt inv DVDD OUT IN DGND
*.PININFO DVDD:B DGND:B OUT:O IN:I
XM1 OUT IN DVDD DVDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.84 nf=1 m=1
XM2 OUT IN DGND DGND sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 m=1
.ends
.end
