** sch_path: /home/ee24s053/ee5311-2025/tut6/sim/pre_layout/fa.sch
.subckt fa DVDD a b cin sum_n cout_n DGND
*.PININFO DVDD:B DGND:B sum_n:O cout_n:O a:I b:I cin:I
XM3 net5 a DGND DGND sky130_fd_pr__nfet_01v8 L=0.15 W=1.68 nf=1 m=1
XM7 cout_n cin net5 DGND sky130_fd_pr__nfet_01v8 L=0.15 W=0.84 nf=1 m=1
XM8 net5 b DGND DGND sky130_fd_pr__nfet_01v8 L=0.15 W=1.68 nf=1 m=1
XM9 net2 a DGND DGND sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM10 net2 b DGND DGND sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM11 net2 cin DGND DGND sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM12 sum_n cout_n net2 DGND sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM13 sum_n cin net7 DGND sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM14 net7 b net8 DGND sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM15 net8 a DGND DGND sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM16 net3 a DVDD DVDD sky130_fd_pr__pfet_01v8 L=0.15 W=1.68 nf=1 m=1
XM18 net4 a DVDD DVDD sky130_fd_pr__pfet_01v8 L=0.15 W=3.36 nf=1 m=1
XM22 cout_n cin net4 DVDD sky130_fd_pr__pfet_01v8 L=0.15 W=1.68 nf=1 m=1
XM23 net4 b DVDD DVDD sky130_fd_pr__pfet_01v8 L=0.15 W=3.36 nf=1 m=1
XM25 sum_n cin net9 DVDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM26 net9 b net10 DVDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM27 net10 a DVDD DVDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM1 net6 a DGND DGND sky130_fd_pr__nfet_01v8 L=0.15 W=0.84 nf=1 m=1
XM2 cout_n b net3 DVDD sky130_fd_pr__pfet_01v8 L=0.15 W=1.68 nf=1 m=1
XM4 cout_n b net6 DGND sky130_fd_pr__nfet_01v8 L=0.15 W=0.84 nf=1 m=1
XM5 net1 a DVDD DVDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM6 net1 b DVDD DVDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM17 net1 cin DVDD DVDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM19 sum_n cout_n net1 DVDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.42 nf=1 m=1
.ends
.end
