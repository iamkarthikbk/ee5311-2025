* Extracted by KLayout with SKY130 LVS runset on : 28/03/2025 14:08

* cell carry_n
* pin DVDD
* pin cout_n
* pin DGND
* pin a
* pin b
* pin cin
* pin GND
.SUBCKT carry_n DVDD cout_n DGND a b cin GND
* device instance $1 r0 *1 -0.97,0.285 sky130_fd_pr__nfet_01v8
XM$1 DGND a \$I26 GND sky130_fd_pr__nfet_01v8 L=150000 W=840000 AS=252000000000
+ AD=210000000000 PS=2280000 PD=1340000
* device instance $2 r0 *1 -0.32,0.285 sky130_fd_pr__nfet_01v8
XM$2 \$I26 b cout_n GND sky130_fd_pr__nfet_01v8 L=150000 W=840000
+ AS=210000000000 AD=210000000000 PS=1340000 PD=1340000
* device instance $3 r0 *1 0.33,0.285 sky130_fd_pr__nfet_01v8
XM$3 cout_n cin \$7 GND sky130_fd_pr__nfet_01v8 L=150000 W=840000
+ AS=210000000000 AD=210000000000 PS=1340000 PD=1340000
* device instance $4 r0 *1 0.98,0.285 sky130_fd_pr__nfet_01v8
XM$4 \$7 b DGND GND sky130_fd_pr__nfet_01v8 L=150000 W=1680000 AS=420000000000
+ AD=420000000000 PS=2680000 PD=2680000
* device instance $6 r0 *1 2.28,0.285 sky130_fd_pr__nfet_01v8
XM$6 \$7 a DGND GND sky130_fd_pr__nfet_01v8 L=150000 W=1680000 AS=420000000000
+ AD=462000000000 PS=2680000 PD=3620000
* device instance $8 r0 *1 -0.97,1.755 sky130_fd_pr__pfet_01v8
XM$8 DVDD a \$5 DVDD sky130_fd_pr__pfet_01v8 L=150000 W=1680000 AS=462000000000
+ AD=462000000000 PS=3620000 PD=3620000
* device instance $9 r0 *1 -0.32,1.755 sky130_fd_pr__pfet_01v8
XM$9 \$5 b cout_n DVDD sky130_fd_pr__pfet_01v8 L=150000 W=1680000
+ AS=420000000000 AD=420000000000 PS=2680000 PD=2680000
* device instance $10 r0 *1 0.33,1.755 sky130_fd_pr__pfet_01v8
XM$10 cout_n cin \$2 DVDD sky130_fd_pr__pfet_01v8 L=150000 W=1680000
+ AS=420000000000 AD=420000000000 PS=2680000 PD=2680000
* device instance $11 r0 *1 0.98,1.755 sky130_fd_pr__pfet_01v8
XM$11 \$2 b DVDD DVDD sky130_fd_pr__pfet_01v8 L=150000 W=3360000
+ AS=840000000000 AD=840000000000 PS=5360000 PD=5360000
* device instance $13 r0 *1 2.28,1.755 sky130_fd_pr__pfet_01v8
XM$13 \$2 a DVDD DVDD sky130_fd_pr__pfet_01v8 L=150000 W=1680000
+ AS=420000000000 AD=420000000000 PS=2680000 PD=2680000
* device instance $15 r0 *1 3.58,1.755 sky130_fd_pr__pfet_01v8
XM$15 \$2 a \$I27 DVDD sky130_fd_pr__pfet_01v8 L=150000 W=1680000
+ AS=420000000000 AD=420000000000 PS=2680000 PD=2680000
.ENDS carry_n
