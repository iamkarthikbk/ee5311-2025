* NGSPICE file created from nand2x1.ext - technology: sky130A

.subckt nand2x1 DGND DVDD B A F
X0 F A a_n694_n141# DGND sky130_fd_pr__nfet_01v8 ad=0.21 pd=1.34 as=0.252 ps=2.28 w=0.84 l=0.15
X1 a_n694_n141# A F DGND sky130_fd_pr__nfet_01v8 ad=0.252 pd=2.28 as=0.21 ps=1.34 w=0.84 l=0.15
X2 F A DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.21 pd=1.34 as=0.252 ps=2.28 w=0.84 l=0.15
X3 DVDD A F DVDD sky130_fd_pr__pfet_01v8 ad=0.5166 pd=2.07 as=0.21 ps=1.34 w=0.84 l=0.15
X4 a_n694_n141# B DGND DGND sky130_fd_pr__nfet_01v8 ad=0.21 pd=1.34 as=0.252 ps=2.28 w=0.84 l=0.15
X5 F B DVDD DVDD sky130_fd_pr__pfet_01v8 ad=0.21 pd=1.34 as=0.5166 ps=2.07 w=0.84 l=0.15
X6 DGND B a_n694_n141# DGND sky130_fd_pr__nfet_01v8 ad=0.252 pd=2.28 as=0.21 ps=1.34 w=0.84 l=0.15
X7 DVDD B F DVDD sky130_fd_pr__pfet_01v8 ad=0.252 pd=2.28 as=0.21 ps=1.34 w=0.84 l=0.15
.ends

