** sch_path: /home/ee24s053/ee5311-2025/tut6/rca/incr/rca8b.sch
.subckt rca8b cin a1 b1 DVDD DGND s1 a2 b2 s2 a3 b3 s3 a4 b4 s4 a5 b5 s5 a6 b6 s6 a7 b7 s7 cout a8 b8 s8
*.PININFO cin:I a1:I b1:I DVDD:B DGND:B s1:O a2:I b2:I s2:O a3:I b3:I s3:O a4:I b4:I s4:O a5:I b5:I s5:O a6:I b6:I s6:O a7:I b7:I
*+ s7:O cout:O a8:I b8:I s8:O
x2 DVDD a1 b1 net1 cin DGND carry_n
x4 DVDD a1 b1 s1 cin net1 DGND sum_n
x1 DVDD a2 net3 DGND invx1
x3 DVDD a2 net2 DGND invx1
x5 DVDD b2 net4 DGND invx1
x6 DVDD b2 net5 DGND invx1
x7 DVDD net2 net4 net6 net1 DGND carry_n
x8 DVDD net3 net5 s2 net1 net6 DGND sum_n
x9 DVDD a3 b3 net7 net6 DGND carry_n
x10 DVDD a3 b3 s3 net6 net7 DGND sum_n
x11 DVDD a4 net9 DGND invx1
x12 DVDD a4 net8 DGND invx1
x13 DVDD b4 net10 DGND invx1
x14 DVDD b4 net11 DGND invx1
x15 DVDD net8 net10 net12 net7 DGND carry_n
x16 DVDD net9 net11 s4 net7 net12 DGND sum_n
x17 DVDD a5 b5 net13 net12 DGND carry_n
x18 DVDD a5 b5 s5 net12 net13 DGND sum_n
x19 DVDD a6 net15 DGND invx1
x20 DVDD a6 net14 DGND invx1
x21 DVDD b6 net16 DGND invx1
x22 DVDD b6 net17 DGND invx1
x23 DVDD net14 net16 net18 net13 DGND carry_n
x24 DVDD net15 net17 s6 net13 net18 DGND sum_n
x25 DVDD a7 b7 net19 net18 DGND carry_n
x26 DVDD a7 b7 s7 net18 net19 DGND sum_n
x27 DVDD a8 net21 DGND invx1
x28 DVDD a8 net20 DGND invx1
x29 DVDD b8 net22 DGND invx1
x30 DVDD b8 net23 DGND invx1
x31 DVDD net20 net22 cout net19 DGND carry_n
x32 DVDD net21 net23 s8 net19 cout DGND sum_n
.ends

* expanding   symbol:  carry_n.sym # of pins=6
** sym_path: /home/ee24s053/ee5311-2025/tut6/rca/incr/carry_n.sym
** sch_path: /home/ee24s053/ee5311-2025/tut6/rca/incr/carry_n.sch
.subckt carry_n DVDD a b cout_n cin DGND
*.PININFO a:I b:I cin:I DGND:B DVDD:B cout_n:O
XM1 net4 a DVDD DVDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM2 net4 a DVDD DVDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM3 net3 a DVDD DVDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM4 net3 a DVDD DVDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM11 cout_n b net4 DVDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM12 cout_n b net4 DVDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM13 cout_n cin net3 DVDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM14 cout_n cin net3 DVDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM25 cout_n b net1 DGND sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM26 net1 a DGND DGND sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM27 cout_n cin net2 DGND sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM28 net2 a DGND DGND sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM5 net3 a DVDD DVDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM6 net3 a DVDD DVDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM7 net3 b DVDD DVDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM8 net3 b DVDD DVDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM9 net3 b DVDD DVDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM10 net3 b DVDD DVDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM29 net2 a DGND DGND sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM30 net2 b DGND DGND sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM31 net2 b DGND DGND sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 m=1
.ends


* expanding   symbol:  sum_n.sym # of pins=7
** sym_path: /home/ee24s053/ee5311-2025/tut6/rca/incr/sum_n.sym
** sch_path: /home/ee24s053/ee5311-2025/tut6/rca/incr/sum_n.sch
.subckt sum_n DVDD a b sum_n cin cout_in DGND
*.PININFO a:I b:I cin:I DGND:B cout_in:I DVDD:B sum_n:O
XM1 net1 a DGND DGND sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM2 net1 b DGND DGND sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM3 net1 cin DGND DGND sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM4 net3 a DGND DGND sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM5 net2 b net3 DGND sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM6 sum_n cin net2 DGND sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM7 sum_n cout_in net1 DGND sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM8 sum_n cout_in net4 DVDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM9 sum_n cin net6 DVDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM10 net6 b net5 DVDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM11 net5 a DVDD DVDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM12 net4 cin DVDD DVDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM13 net4 b DVDD DVDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM14 net4 a DVDD DVDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.42 nf=1 m=1
.ends


* expanding   symbol:  invx1.sym # of pins=4
** sym_path: /home/ee24s053/ee5311-2025/tut6/rca/incr/invx1.sym
** sch_path: /home/ee24s053/ee5311-2025/tut6/rca/incr/invx1.sch
.subckt invx1 DVDD in out DGND
*.PININFO in:I out:O DVDD:B DGND:B
XM2 out in DVDD DVDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.84 nf=1 m=1
XM1 out in DGND DGND sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 m=1
.ends

.end
