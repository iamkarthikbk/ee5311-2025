* NGSPICE file created from ro7.ext - technology: sky130A
.subckt ro7 DVDD vout DGND
X0 a_n1524_n46# a_n1822_n46# DGND.t13 DGND.t12 sky130_fd_pr__nfet_01v8 ad=0.126 pd=1.44 as=0.126 ps=1.44 w=0.42 l=0.15
X1 a_n332_n46# a_n630_n46# DGND.t9 DGND.t8 sky130_fd_pr__nfet_01v8 ad=0.126 pd=1.44 as=0.126 ps=1.44 w=0.42 l=0.15
X2 a_n928_n46# a_n1226_n46# DVDD.t9 DVDD.t8 sky130_fd_pr__pfet_01v8 ad=0.252 pd=2.28 as=0.252 ps=2.28 w=0.84 l=0.15
X3 vout.t1 a_n332_n46# DGND.t3 DGND.t2 sky130_fd_pr__nfet_01v8 ad=0.126 pd=1.44 as=0.126 ps=1.44 w=0.42 l=0.15
X4 a_n1226_n46# a_n1524_n46# DGND.t1 DGND.t0 sky130_fd_pr__nfet_01v8 ad=0.126 pd=1.44 as=0.126 ps=1.44 w=0.42 l=0.15
X5 a_n1822_n46# vout.t2 DVDD.t7 DVDD.t6 sky130_fd_pr__pfet_01v8 ad=0.252 pd=2.28 as=0.252 ps=2.28 w=0.84 l=0.15
X6 a_n630_n46# a_n928_n46# DVDD.t5 DVDD.t4 sky130_fd_pr__pfet_01v8 ad=0.252 pd=2.28 as=0.252 ps=2.28 w=0.84 l=0.15
X7 a_n1524_n46# a_n1822_n46# DVDD.t13 DVDD.t12 sky130_fd_pr__pfet_01v8 ad=0.252 pd=2.28 as=0.252 ps=2.28 w=0.84 l=0.15
X8 a_n928_n46# a_n1226_n46# DGND.t7 DGND.t6 sky130_fd_pr__nfet_01v8 ad=0.126 pd=1.44 as=0.126 ps=1.44 w=0.42 l=0.15
X9 a_n332_n46# a_n630_n46# DVDD.t11 DVDD.t10 sky130_fd_pr__pfet_01v8 ad=0.252 pd=2.28 as=0.252 ps=2.28 w=0.84 l=0.15
X10 vout.t0 a_n332_n46# DVDD.t3 DVDD.t2 sky130_fd_pr__pfet_01v8 ad=0.252 pd=2.28 as=0.252 ps=2.28 w=0.84 l=0.15
X11 a_n1822_n46# vout.t3 DGND.t11 DGND.t10 sky130_fd_pr__nfet_01v8 ad=0.126 pd=1.44 as=0.126 ps=1.44 w=0.42 l=0.15
X12 a_n1226_n46# a_n1524_n46# DVDD.t1 DVDD.t0 sky130_fd_pr__pfet_01v8 ad=0.252 pd=2.28 as=0.252 ps=2.28 w=0.84 l=0.15
X13 a_n630_n46# a_n928_n46# DGND.t5 DGND.t4 sky130_fd_pr__nfet_01v8 ad=0.126 pd=1.44 as=0.126 ps=1.44 w=0.42 l=0.15
R0 DGND.n6 DGND.t2 4667.36
R1 DGND.t2 DGND.t8 4284.97
R2 DGND.t8 DGND.t4 4284.97
R3 DGND.t4 DGND.t6 4284.97
R4 DGND.t6 DGND.t0 4284.97
R5 DGND.t0 DGND.t12 4284.97
R6 DGND.t12 DGND.t10 4284.97
R7 DGND.n0 DGND.t11 282.904
R8 DGND.n0 DGND.t13 282.515
R9 DGND.n1 DGND.t1 282.515
R10 DGND.n2 DGND.t7 282.515
R11 DGND.n3 DGND.t5 282.515
R12 DGND.n4 DGND.t9 282.515
R13 DGND.n5 DGND.t3 282.515
R14 DGND.n5 DGND.n4 0.388521
R15 DGND.n4 DGND.n3 0.388521
R16 DGND.n3 DGND.n2 0.388521
R17 DGND.n2 DGND.n1 0.388521
R18 DGND.n1 DGND.n0 0.388521
R19 DGND.n6 DGND.n5 0.371594
R20 DGND DGND.n6 0.00180208
R21 DVDD DVDD.t2 945.404
R22 DVDD.t2 DVDD.t10 873.765
R23 DVDD.t10 DVDD.t4 873.765
R24 DVDD.t4 DVDD.t8 873.765
R25 DVDD.t8 DVDD.t0 873.765
R26 DVDD.t0 DVDD.t12 873.765
R27 DVDD.t12 DVDD.t6 873.765
R28 DVDD.n0 DVDD.t7 406.897
R29 DVDD.n0 DVDD.t13 406.509
R30 DVDD.n1 DVDD.t1 406.509
R31 DVDD.n2 DVDD.t9 406.509
R32 DVDD.n3 DVDD.t5 406.509
R33 DVDD.n4 DVDD.t11 406.509
R34 DVDD.n5 DVDD.t3 406.509
R35 DVDD.n5 DVDD.n4 0.388521
R36 DVDD.n4 DVDD.n3 0.388521
R37 DVDD.n3 DVDD.n2 0.388521
R38 DVDD.n2 DVDD.n1 0.388521
R39 DVDD.n1 DVDD.n0 0.388521
R40 DVDD DVDD.n5 0.370292
R41 vout.n2 vout.t0 414.344
R42 vout.n0 vout.t2 303.99
R43 vout.n2 vout.t1 259.481
R44 vout.n4 vout.n0 166.407
R45 vout.n0 vout.t3 144.929
R46 vout.n3 vout.n2 12.8005
R47 vout.n4 vout.n3 9.3005
R48 vout.n3 vout.n1 0.557022
R49 vout vout.n4 0.00593478
C0 a_n928_n46# DVDD 0.221672f
C1 a_n630_n46# a_n928_n46# 0.072255f
C2 vout a_n928_n46# 0.064931f
C3 a_n1226_n46# a_n928_n46# 0.072255f
C4 a_n1822_n46# DVDD 0.219036f
C5 a_n1524_n46# a_n1822_n46# 0.072255f
C6 a_n1822_n46# vout 0.12314f
C7 DVDD a_n332_n46# 0.22299f
C8 a_n630_n46# DVDD 0.221672f
C9 a_n1524_n46# DVDD 0.221672f
C10 vout DVDD 0.592581f
C11 a_n630_n46# a_n332_n46# 0.072255f
C12 vout a_n332_n46# 0.119328f
C13 a_n630_n46# vout 0.064931f
C14 a_n1524_n46# vout 0.064931f
C15 a_n1226_n46# DVDD 0.221672f
C16 a_n1524_n46# a_n1226_n46# 0.072255f
C17 vout a_n1226_n46# 0.064931f
C18 vout DGND 0.920549f
C19 DVDD DGND 2.91043f
C20 a_n332_n46# DGND 0.34096f
C21 a_n630_n46# DGND 0.324985f
C22 a_n928_n46# DGND 0.324985f
C23 a_n1226_n46# DGND 0.324985f
C24 a_n1524_n46# DGND 0.324985f
C25 a_n1822_n46# DGND 0.344123f
.ends
