** sch_path: /home/ee24s053/ee5311-2025/tut6/again/sum/sum.sch
.subckt sum an bn cin DGND cout_in DVDD sum_n
*.PININFO an:I bn:I cin:I DGND:B cout_in:I DVDD:B sum_n:O
XM1 net1 a DGND DGND sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM2 net1 b DGND DGND sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM3 net1 cin DGND DGND sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM4 net3 a DGND DGND sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM5 net2 b net3 DGND sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM6 sum_n cin net2 DGND sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM7 sum_n cout_in net1 DGND sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM8 sum_n cout_in net4 DVDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 m=1
XM9 sum_n cin net6 DVDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 m=1
XM10 net6 b net5 DVDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 m=1
XM11 net5 a DVDD DVDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 m=1
XM12 net4 cin DVDD DVDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 m=1
XM13 net4 b DVDD DVDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 m=1
XM14 net4 a DVDD DVDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 m=1
XM15 a an DVDD DVDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 m=1
XM16 a an DGND DGND sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM17 b bn DVDD DVDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 m=1
XM18 b bn DGND DGND sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 m=1
.ends
.end
