** sch_path: /home/ee24s053/ee5311-2025/tut5/inv/sim/post-layout/delay.sch
**.subckt delay inp outp del

x1 VDD vout vin GND inv_nosubckt
x2 VDD net1 vout GND inv_nosubckt
V1 vin GND PULSE(0 1.8 10ps 5ps 5ps 100ps 250ps)
V2 VDD GND 1.8
**** begin user architecture code
.lib /cad/share/pdk/sky130B/libs.tech/combined/sky130.lib.spice tt


.include /home/ee24s053/ee5311-2025/tut5/inv/prim/inv_extracted.spice
.control
tran 0.01p 250p
plot v(vout) v(vin)
meas tran thl trig v(vin) val=0.9 rise=1 targ v(vout) val=0.9 fall=1
meas tran tlh trig v(vin) val=0.9 fall=1 targ v(vout) val=0.9 rise=1
let delay = ($&tlh + $&thl) /2
echo delay: $&delay
.endc


**** end user architecture code
**.ends
.GLOBAL VDD
.GLOBAL GND
.end
