** sch_path: /home/ee24s053/ee5311-2025/tut6/again/sim/adder_parasitics.sch
**.subckt adder_parasitics
x1 VDD a_tap b_tap cout_n_tap cin_tap GND carry_n
x2 VDD a_tap b_tap sum_n_tap cin_tap cout_n_tap GND sum_n
x3 VDD net2 net3 net1 cout_n_tap GND carry
x4 VDD net2 net4 net3 cout_n_tap net1 GND sum
V1 a_tap GND 0
V2 b_tap GND 1.8
V3 cin_tap GND PULSE(0 1.8 0 50ns 50ns 1us 2us)
V4 net2 GND 0
V5 net3 GND 1.8
V6 VDD GND 1.8
**** begin user architecture code


.include /home/ee24s053/ee5311-2025/tut6/again/sum/sum_extracted.spice
.include /home/ee24s053/ee5311-2025/tut6/again/sum_n/sum_n_extracted.spice
.include /home/ee24s053/ee5311-2025/tut6/again/carry/carry_extracted.spice
.include /home/ee24s053/ee5311-2025/tut6/again/carry_n/carry_n_extracted.spice
.control
tran 1n 20u
plot v(a_tap) v(b_tap) v(cin_tap)
plot v(sum_n_tap) v(cout_n_tap)
meas tran tlh_carry trig v(cin_tap) val=0.9 rise=1 targ v(cout_n_tap) val=0.9 rise=1
meas tran thl_carry trig v(cin_tap) val=0.9 fall=1 targ v(cout_n_tap) val=0.9 fall=1
let carry_delay = ($&tlh_carry + $&thl_carry)/2
echo carry delay: $&carry_delay
meas tran tlh_sum trig v(cin_tap) val=0.9 rise=1 targ v(sum_n_tap) val=0.9 rise=1
meas tran thl_sum trig v(cin_tap) val=0.9 fall=1 targ v(sum_n_tap) val=0.9 fall=1
let sum_delay = ($&tlh_sum + $&thl_sum)/2
echo sum delay: $&sum_delay
.endc

.lib /cad/share/pdk/sky130B/libs.tech/combined/sky130.lib.spice tt
**** end user architecture code
**.ends
.GLOBAL VDD
.GLOBAL GND
.end
