** sch_path: /home/ee24s053/ee5311-2025/tut1/pmos/expt2/expt2.sch
**.subckt expt2
Vin1 Vin GND 1.8
Vdd1 net1 GND 1.8
XM1 GND Vin net1 VDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
**** begin user architecture code
.lib /cad/share/pdk/sky130B/libs.tech/combined/sky130.lib.spice tt

.control
let Vgs=0.6
repeat 4
  alter Vin1 $&Vgs
  dc Vdd1 0 1.8 0.02
  let Vgs=Vgs+0.4
end
plot dc1.I(Vdd1)*-1 dc2.I(Vdd1)*-1 dc3.I(Vdd1)*-1 dc4.I(Vdd1)*-1
set filetype=ascii
wrdata pmos_ids_vds.txt dc1.I(Vdd1)*-1 dc2.I(Vdd1)*-1 dc3.I(Vdd1)*-1 dc4.I(Vdd1)*-1
.endc

**** end user architecture code
**.ends
.GLOBAL GND
.end
