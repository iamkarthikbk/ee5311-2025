** sch_path: /home/ee24s053/ee5311-2025/tut5/ro7/cell/ro7.sch
.subckt ro7

Vdd1 VDD GND {vdd_val}
x1 VDD net1 vout GND inv
x2 VDD net2 net1 GND inv
x3 VDD net3 net2 GND inv
x4 VDD net4 net3 GND inv
x5 VDD net5 net4 GND inv
x6 VDD net6 net5 GND inv
x7 VDD vout net6 GND inv
**** begin user architecture code
.lib /cad/share/pdk/sky130B/libs.tech/combined/sky130.lib.spice tt


.param vdd_val = 1.8
.ic v(vout) = 0
.control
let lv_iters = 9
let v_vdd = vector(lv_iters)
let v_period = vector(lv_iters)
let v_freq = vector(lv_iters)
let lv_index = 0
while lv_index < lv_iters
	let lv_vdd = 1.0 + (lv_index * 0.1)
	let vhalf = lv_vdd / 2
	alterparam vdd_val = $&lv_vdd
	reset
	tran 1p 10n
	meas tran prd trig v(vout) val=vhalf rise=3 targ v(vout) val=vhalf rise=4
	let v_period[lv_index] = $&prd
	let v_freq[lv_index] = 1/$&prd
	let v_vdd[lv_index] = $&lv_vdd
	let lv_index = lv_index + 1
end
plot v_period vs v_vdd
plot v_freq vs v_vdd
.endc


**** end user architecture code
.ends

* expanding   symbol:  /home/ee24s053/ee5311-2025/tut5/inv/cell/subcircuit/inv.sym # of pins=4
** sym_path: /home/ee24s053/ee5311-2025/tut5/inv/cell/subcircuit/inv.sym
** sch_path: /home/ee24s053/ee5311-2025/tut5/inv/cell/subcircuit/inv.sch
.subckt inv DVDD OUT IN DGND
*.PININFO DVDD:B DGND:B OUT:O IN:I
XM1 OUT IN DVDD DVDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.84 nf=1 m=1
XM2 OUT IN DGND DGND sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 m=1
.ends

.GLOBAL VDD
.GLOBAL GND
.end
