* NGSPICE file created from nand2x1.ext - technology: sky130A

.subckt pfet a_90_0# a_60_n40# w_n63_n78# a_220_0# a_0_0# a_190_n40#
X0 a_90_0# a_60_n40# a_0_0# w_n63_n78# sky130_fd_pr__pfet_01v8 ad=0.21 pd=1.34 as=0.252 ps=2.28 w=0.84 l=0.15
X1 a_220_0# a_190_n40# a_90_0# w_n63_n78# sky130_fd_pr__pfet_01v8 ad=0.252 pd=2.28 as=0.21 ps=1.34 w=0.84 l=0.15
.ends

.subckt nfet a_90_0# a_60_n40# a_220_0# a_0_0# a_190_n40# VSUBS
X0 a_90_0# a_60_n40# a_0_0# VSUBS sky130_fd_pr__nfet_01v8 ad=0.21 pd=1.34 as=0.252 ps=2.28 w=0.84 l=0.15
X1 a_220_0# a_190_n40# a_90_0# VSUBS sky130_fd_pr__nfet_01v8 ad=0.252 pd=2.28 as=0.21 ps=1.34 w=0.84 l=0.15
.ends

.subckt nand2x1 DGND DVDD B A F
Xpfet_0 F A DVDD DVDD DVDD A pfet
Xpfet_1 F B DVDD DVDD DVDD B pfet
Xnfet_0 F A DGND DGND A DGND nfet
Xnfet_1 DGND B DGND DGND B DGND nfet
.ends

