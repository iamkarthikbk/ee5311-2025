** sch_path: /home/ee24s053/ee5311-2025/tut2/expt2_1/expt2_1.sch
**.subckt expt2_1
XM1 Vout Vin GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
Vin1 Vin GND 1.8
XM2 Vout Vin VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
Vdd1 VDD GND 1.8
**** begin user architecture code
.lib /cad/share/pdk/sky130B/libs.tech/combined/sky130.lib.spice tt

.control
let vds = 0.2
set cache = ''
let index = 1
let N = 10
let imax = vector(N)
while index le N
  alter Vdd1 $&vds
  dc Vin1 0 $&vds 0.01
  set cache = ( $cache dc($&index) .v(Vout) )
  let imax[index - 1] = abs(vecmin(dc{$&index}.i(Vdd1)))
  let vds = vds + 0.2
  let index = index + 1
end
plot $cache
.endc

**** end user architecture code
**.ends
.GLOBAL GND
.end
