* NGSPICE file created from invx1.ext - technology: sky130A
.subckt invx1 in out DVDD DGND
X0 out.t0 in.t0 DGND.t1 DGND.t0 sky130_fd_pr__nfet_01v8 ad=0.126 pd=1.44 as=0.126 ps=1.44 w=0.42 l=0.15
X1 out.t1 in.t1 DVDD.t1 DVDD.t0 sky130_fd_pr__pfet_01v8 ad=0.252 pd=2.28 as=0.252 ps=2.28 w=0.84 l=0.15
R0 in.n0 in.t1 240.096
R1 in.n0 in.t0 175.831
R2 in in.n0 152.948
R3 DGND DGND.t0 4921.89
R4 DGND DGND.t1 272.351
R5 out.t1 out 705.836
R6 out.n1 out.t1 703.201
R7 out.n0 out.t0 227.857
R8 out out.n1 6.4005
R9 out.n0 out 6.4005
R10 out.n1 out 1.12991
R11 out out.n0 1.12991
R12 DVDD DVDD.t1 405.103
R13 DVDD DVDD.t0 274.622
C0 out DVDD 0.072397f
C1 in DVDD 0.106979f
C2 in out 0.036249f
C3 out DGND 0.144607f
C4 in DGND 0.226044f
C5 DVDD DGND 0.756609f
.ends
