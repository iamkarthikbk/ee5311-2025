** sch_path: /home/ee24s053/ee5311-2025/mywork/nor2x1/nor2x1.sch
.subckt nor2x1 DVDD DGND A F B
*.PININFO DVDD:B DGND:B A:I F:O B:I
XM1 net1 A DVDD DVDD sky130_fd_pr__pfet_01v8 L=0.15 W=1.68 nf=4 m=1
XM2 F B net1 DVDD sky130_fd_pr__pfet_01v8 L=0.15 W=1.68 nf=4 m=1
XM3 F A DGND DGND sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 m=1
XM4 F B DGND DGND sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 m=1
.ends
.end
