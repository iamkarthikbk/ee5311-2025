** sch_path: /home/ee24s053/ee5311-2025/tut6/sim/pre_layout/incr/msym-fa-sum-pdn.sch
.subckt msym-fa-sum-pdn out a b c1 c2 bot
*.PININFO out:O a:I b:I c1:I c2:I bot:B
XM1 net1 c1 bot bot sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM2 net1 b bot bot sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM3 net1 a bot bot sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM4 out c2 net1 bot sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM5 net2 a bot bot sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM6 net3 b net2 bot sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM7 out c1 net3 bot sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM8 out c2 net6 net4 sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 m=1
XM9 net6 a net4 net4 sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 m=1
XM10 net6 b net4 net4 sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 m=1
XM11 net6 c1 net4 net4 sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 m=1
XM12 net5 a net4 net4 sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 m=1
XM13 net7 b net5 net4 sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 m=1
XM14 out c1 net7 net4 sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 m=1
.ends
.end
