* NGSPICE file created from inv.ext - technology: sky130A

.subckt pfet$1 a_90_0# a_60_n40# w_n63_n78# a_0_0#
X0 a_90_0# a_60_n40# a_0_0# w_n63_n78# sky130_fd_pr__pfet_01v8 ad=0.252 pd=2.28 as=0.252 ps=2.28 w=0.84 l=0.15
.ends

.subckt inv IN OUT DVDD DGND
Xpfet$1_0 OUT IN DVDD DVDD pfet$1
X0 OUT IN DGND DGND sky130_fd_pr__nfet_01v8 ad=0.126 pd=1.44 as=0.126 ps=1.44 w=0.42 l=0.15
.ends

