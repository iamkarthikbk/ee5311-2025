** sch_path: /home/ee24s053/ee5311-2025/tut1/pmos/expt1_0/expt1_0.sch
**.subckt expt1_0
Vin1 Vin GND 0
XM1 Vin Vin GND VDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
**** begin user architecture code
.lib /cad/share/pdk/sky130B/libs.tech/combined/sky130.lib.spice tt

.control
set filetype=ascii
dc Vin1 0 -1.8 -0.01
wrdata pmos_ids_vgs.txt -I(Vin1)
.endc

**** end user architecture code
**.ends
.GLOBAL GND
.end
