* NGSPICE file created from ro7.ext - technology: sky130A

.subckt pfet$1 a_90_0# a_60_n40# w_n63_n78# a_0_0#
X0 a_90_0# a_60_n40# a_0_0# w_n63_n78# sky130_fd_pr__pfet_01v8 ad=0.252 pd=2.28 as=0.252 ps=2.28 w=0.84 l=0.15
.ends

.subckt inv_wo_tap OUT pfet$1_0/w_n63_n78# DVDD DGND IN VSUBS
Xpfet$1_0 OUT IN pfet$1_0/w_n63_n78# DVDD pfet$1
X0 OUT IN DGND VSUBS sky130_fd_pr__nfet_01v8 ad=0.126 pd=1.44 as=0.126 ps=1.44 w=0.42 l=0.15
.ends

.subckt ro7 vout DVDD DGND
Xinv_wo_tap_0 inv_wo_tap_1/IN DVDD DVDD DGND vout DGND inv_wo_tap
Xinv_wo_tap_1 inv_wo_tap_2/IN DVDD DVDD DGND inv_wo_tap_1/IN DGND inv_wo_tap
Xinv_wo_tap_2 inv_wo_tap_3/IN DVDD DVDD DGND inv_wo_tap_2/IN DGND inv_wo_tap
Xinv_wo_tap_4 inv_wo_tap_5/IN DVDD DVDD DGND inv_wo_tap_4/IN DGND inv_wo_tap
Xinv_wo_tap_3 inv_wo_tap_4/IN DVDD DVDD DGND inv_wo_tap_3/IN DGND inv_wo_tap
Xinv_wo_tap_5 inv_wo_tap_6/IN DVDD DVDD DGND inv_wo_tap_5/IN DGND inv_wo_tap
Xinv_wo_tap_6 vout DVDD DVDD DGND inv_wo_tap_6/IN DGND inv_wo_tap
.ends

